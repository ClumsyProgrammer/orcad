** Profile: "ROOT-vdd_sweep"  [ C:\Users\katerina\Desktop\synodeutiko_yliko\gates\ccdd\XOR\45nm\ccdd_xor_45-pspicefiles\root\vdd_sweep.sim ] 

** Creating circuit file "vdd_sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Users/katerina/Desktop/ptyxiaki/ptm_library/PTM_Models.lib" 
.STMLIB "../../../ccdd_xor_45-pspicefiles/ccdd_xor_45.stl" 
* From [PSPICE NETLIST] section of C:\Users\katerina\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1.2ns 0 
.STEP LIN PARAM vdd_nominal 1 2.5 0.5 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\ROOT.net" 


.END
