** Profile: "GATE-gate"  [ C:\Users\katerina\Desktop\synodeutiko_yliko\gates\dcml\XOR\45nm\dcml_xor_45-pspicefiles\gate\gate.sim ] 

** Creating circuit file "gate.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Users/katerina/Desktop/ptyxiaki/ptm_library/PTM_Models.lib" 
.STMLIB "../../../dcml_xor_45-pspicefiles/dcml_xor_45.stl" 
* From [PSPICE NETLIST] section of C:\Users\katerina\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\GATE.net" 


.END
